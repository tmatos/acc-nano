// ----------------------------------------------------------------------------
// LegUp High-Level Synthesis Tool Version 7.2 (http://legupcomputing.com)
// Copyright (c) 2015-2019 LegUp Computing Inc. All Rights Reserved.
// For technical issues, please contact: support@legupcomputing.com
// For general inquiries, please contact: info@legupcomputing.com
// Date: Mon Aug 12 04:54:19 2019
// ----------------------------------------------------------------------------

`define MEMORY_CONTROLLER_ADDR_SIZE 32

// This directory contains the memory initialization files generated by LegUp.
// This relative path is used by ModelSim and FPGA synthesis tool.
`define MEM_INIT_DIR "../mem_init/"

`timescale 1 ns / 1 ns

module kernel_atax_top
(
	clk,
	reset,
	start,
	finish,
	main_y_write_enable_a,
	main_y_in_a,
	main_y_byteena_a,
	main_y_enable_a,
	main_y_address_a,
	main_y_out_a,
	main_y_write_enable_b,
	main_y_in_b,
	main_y_byteena_b,
	main_y_enable_b,
	main_y_address_b,
	main_y_out_b,
	main_x_write_enable_a,
	main_x_in_a,
	main_x_byteena_a,
	main_x_enable_a,
	main_x_address_a,
	main_x_out_a,
	main_x_write_enable_b,
	main_x_in_b,
	main_x_byteena_b,
	main_x_enable_b,
	main_x_address_b,
	main_x_out_b,
	main_A_a0_a0_write_enable_a,
	main_A_a0_a0_in_a,
	main_A_a0_a0_byteena_a,
	main_A_a0_a0_enable_a,
	main_A_a0_a0_address_a,
	main_A_a0_a0_out_a,
	main_A_a0_a0_write_enable_b,
	main_A_a0_a0_in_b,
	main_A_a0_a0_byteena_b,
	main_A_a0_a0_enable_b,
	main_A_a0_a0_address_b,
	main_A_a0_a0_out_b
);

input  clk;
input  reset;
input  start;
output reg  finish;
output reg  main_y_write_enable_a;
output reg [63:0] main_y_in_a;
output reg  main_y_byteena_a;
output  main_y_enable_a;
output reg [4:0] main_y_address_a;
input [63:0] main_y_out_a;
output reg  main_y_write_enable_b;
output reg [63:0] main_y_in_b;
output reg  main_y_byteena_b;
output  main_y_enable_b;
output reg [4:0] main_y_address_b;
input [63:0] main_y_out_b;
output reg  main_x_write_enable_a;
output reg [63:0] main_x_in_a;
output reg  main_x_byteena_a;
output  main_x_enable_a;
output reg [4:0] main_x_address_a;
input [63:0] main_x_out_a;
output reg  main_x_write_enable_b;
output reg [63:0] main_x_in_b;
output reg  main_x_byteena_b;
output  main_x_enable_b;
output reg [4:0] main_x_address_b;
input [63:0] main_x_out_b;
output reg  main_A_a0_a0_write_enable_a;
output reg [63:0] main_A_a0_a0_in_a;
output reg  main_A_a0_a0_byteena_a;
output  main_A_a0_a0_enable_a;
output reg [9:0] main_A_a0_a0_address_a;
input [63:0] main_A_a0_a0_out_a;
output reg  main_A_a0_a0_write_enable_b;
output reg [63:0] main_A_a0_a0_in_b;
output reg  main_A_a0_a0_byteena_b;
output  main_A_a0_a0_enable_b;
output reg [9:0] main_A_a0_a0_address_b;
input [63:0] main_A_a0_a0_out_b;
reg  kernel_atax_inst_clk;
reg  kernel_atax_inst_reset;
reg  kernel_atax_inst_start;
wire  kernel_atax_inst_finish;
wire  kernel_atax_inst_main_y_write_enable_a;
wire [63:0] kernel_atax_inst_main_y_in_a;
wire  kernel_atax_inst_main_y_byteena_a;
wire  kernel_atax_inst_main_y_enable_a;
wire [4:0] kernel_atax_inst_main_y_address_a;
reg [63:0] kernel_atax_inst_main_y_out_a;
wire  kernel_atax_inst_main_y_write_enable_b;
wire [63:0] kernel_atax_inst_main_y_in_b;
wire  kernel_atax_inst_main_y_byteena_b;
wire  kernel_atax_inst_main_y_enable_b;
wire [4:0] kernel_atax_inst_main_y_address_b;
reg [63:0] kernel_atax_inst_main_y_out_b;
wire  kernel_atax_inst_main_x_write_enable_a;
wire [63:0] kernel_atax_inst_main_x_in_a;
wire  kernel_atax_inst_main_x_byteena_a;
wire  kernel_atax_inst_main_x_enable_a;
wire [4:0] kernel_atax_inst_main_x_address_a;
reg [63:0] kernel_atax_inst_main_x_out_a;
wire  kernel_atax_inst_main_x_write_enable_b;
wire [63:0] kernel_atax_inst_main_x_in_b;
wire  kernel_atax_inst_main_x_byteena_b;
wire  kernel_atax_inst_main_x_enable_b;
wire [4:0] kernel_atax_inst_main_x_address_b;
reg [63:0] kernel_atax_inst_main_x_out_b;
wire  kernel_atax_inst_main_A_a0_a0_write_enable_a;
wire [63:0] kernel_atax_inst_main_A_a0_a0_in_a;
wire  kernel_atax_inst_main_A_a0_a0_byteena_a;
wire  kernel_atax_inst_main_A_a0_a0_enable_a;
wire [9:0] kernel_atax_inst_main_A_a0_a0_address_a;
reg [63:0] kernel_atax_inst_main_A_a0_a0_out_a;
wire  kernel_atax_inst_main_A_a0_a0_write_enable_b;
wire [63:0] kernel_atax_inst_main_A_a0_a0_in_b;
wire  kernel_atax_inst_main_A_a0_a0_byteena_b;
wire  kernel_atax_inst_main_A_a0_a0_enable_b;
wire [9:0] kernel_atax_inst_main_A_a0_a0_address_b;
reg [63:0] kernel_atax_inst_main_A_a0_a0_out_b;
reg  kernel_atax_inst_finish_reg;


kernel_atax kernel_atax_inst (
	.clk (kernel_atax_inst_clk),
	.reset (kernel_atax_inst_reset),
	.start (kernel_atax_inst_start),
	.finish (kernel_atax_inst_finish),
	.main_y_write_enable_a (kernel_atax_inst_main_y_write_enable_a),
	.main_y_in_a (kernel_atax_inst_main_y_in_a),
	.main_y_byteena_a (kernel_atax_inst_main_y_byteena_a),
	.main_y_enable_a (kernel_atax_inst_main_y_enable_a),
	.main_y_address_a (kernel_atax_inst_main_y_address_a),
	.main_y_out_a (kernel_atax_inst_main_y_out_a),
	.main_y_write_enable_b (kernel_atax_inst_main_y_write_enable_b),
	.main_y_in_b (kernel_atax_inst_main_y_in_b),
	.main_y_byteena_b (kernel_atax_inst_main_y_byteena_b),
	.main_y_enable_b (kernel_atax_inst_main_y_enable_b),
	.main_y_address_b (kernel_atax_inst_main_y_address_b),
	.main_y_out_b (kernel_atax_inst_main_y_out_b),
	.main_x_write_enable_a (kernel_atax_inst_main_x_write_enable_a),
	.main_x_in_a (kernel_atax_inst_main_x_in_a),
	.main_x_byteena_a (kernel_atax_inst_main_x_byteena_a),
	.main_x_enable_a (kernel_atax_inst_main_x_enable_a),
	.main_x_address_a (kernel_atax_inst_main_x_address_a),
	.main_x_out_a (kernel_atax_inst_main_x_out_a),
	.main_x_write_enable_b (kernel_atax_inst_main_x_write_enable_b),
	.main_x_in_b (kernel_atax_inst_main_x_in_b),
	.main_x_byteena_b (kernel_atax_inst_main_x_byteena_b),
	.main_x_enable_b (kernel_atax_inst_main_x_enable_b),
	.main_x_address_b (kernel_atax_inst_main_x_address_b),
	.main_x_out_b (kernel_atax_inst_main_x_out_b),
	.main_A_a0_a0_write_enable_a (kernel_atax_inst_main_A_a0_a0_write_enable_a),
	.main_A_a0_a0_in_a (kernel_atax_inst_main_A_a0_a0_in_a),
	.main_A_a0_a0_byteena_a (kernel_atax_inst_main_A_a0_a0_byteena_a),
	.main_A_a0_a0_enable_a (kernel_atax_inst_main_A_a0_a0_enable_a),
	.main_A_a0_a0_address_a (kernel_atax_inst_main_A_a0_a0_address_a),
	.main_A_a0_a0_out_a (kernel_atax_inst_main_A_a0_a0_out_a),
	.main_A_a0_a0_write_enable_b (kernel_atax_inst_main_A_a0_a0_write_enable_b),
	.main_A_a0_a0_in_b (kernel_atax_inst_main_A_a0_a0_in_b),
	.main_A_a0_a0_byteena_b (kernel_atax_inst_main_A_a0_a0_byteena_b),
	.main_A_a0_a0_enable_b (kernel_atax_inst_main_A_a0_a0_enable_b),
	.main_A_a0_a0_address_b (kernel_atax_inst_main_A_a0_a0_address_b),
	.main_A_a0_a0_out_b (kernel_atax_inst_main_A_a0_a0_out_b)
);



always @(*) begin
	kernel_atax_inst_clk = clk;
end
always @(*) begin
	kernel_atax_inst_reset = reset;
end
always @(*) begin
	kernel_atax_inst_start = start;
end
always @(*) begin
	kernel_atax_inst_main_y_out_a = main_y_out_a;
end
always @(*) begin
	kernel_atax_inst_main_y_out_b = main_y_out_b;
end
always @(*) begin
	kernel_atax_inst_main_x_out_a = main_x_out_a;
end
always @(*) begin
	kernel_atax_inst_main_x_out_b = main_x_out_b;
end
always @(*) begin
	kernel_atax_inst_main_A_a0_a0_out_a = main_A_a0_a0_out_a;
end
always @(*) begin
	kernel_atax_inst_main_A_a0_a0_out_b = main_A_a0_a0_out_b;
end
always @(posedge clk) begin
	if ((reset | kernel_atax_inst_start)) begin
		kernel_atax_inst_finish_reg <= 1'd0;
	end
	if (kernel_atax_inst_finish) begin
		kernel_atax_inst_finish_reg <= 1'd1;
	end
end
always @(*) begin
	finish = kernel_atax_inst_finish;
end
always @(*) begin
	main_y_write_enable_a = kernel_atax_inst_main_y_write_enable_a;
end
always @(*) begin
	main_y_in_a = kernel_atax_inst_main_y_in_a;
end
always @(*) begin
	main_y_byteena_a = kernel_atax_inst_main_y_byteena_a;
end
assign main_y_enable_a = 0;
always @(*) begin
	main_y_address_a = kernel_atax_inst_main_y_address_a;
end
always @(*) begin
	main_y_write_enable_b = kernel_atax_inst_main_y_write_enable_b;
end
always @(*) begin
	main_y_in_b = kernel_atax_inst_main_y_in_b;
end
always @(*) begin
	main_y_byteena_b = kernel_atax_inst_main_y_byteena_b;
end
assign main_y_enable_b = 0;
always @(*) begin
	main_y_address_b = kernel_atax_inst_main_y_address_b;
end
always @(*) begin
	main_x_write_enable_a = kernel_atax_inst_main_x_write_enable_a;
end
always @(*) begin
	main_x_in_a = kernel_atax_inst_main_x_in_a;
end
always @(*) begin
	main_x_byteena_a = kernel_atax_inst_main_x_byteena_a;
end
assign main_x_enable_a = 0;
always @(*) begin
	main_x_address_a = kernel_atax_inst_main_x_address_a;
end
always @(*) begin
	main_x_write_enable_b = kernel_atax_inst_main_x_write_enable_b;
end
always @(*) begin
	main_x_in_b = kernel_atax_inst_main_x_in_b;
end
always @(*) begin
	main_x_byteena_b = kernel_atax_inst_main_x_byteena_b;
end
assign main_x_enable_b = 0;
always @(*) begin
	main_x_address_b = kernel_atax_inst_main_x_address_b;
end
always @(*) begin
	main_A_a0_a0_write_enable_a = kernel_atax_inst_main_A_a0_a0_write_enable_a;
end
always @(*) begin
	main_A_a0_a0_in_a = kernel_atax_inst_main_A_a0_a0_in_a;
end
always @(*) begin
	main_A_a0_a0_byteena_a = kernel_atax_inst_main_A_a0_a0_byteena_a;
end
assign main_A_a0_a0_enable_a = 0;
always @(*) begin
	main_A_a0_a0_address_a = kernel_atax_inst_main_A_a0_a0_address_a;
end
always @(*) begin
	main_A_a0_a0_write_enable_b = kernel_atax_inst_main_A_a0_a0_write_enable_b;
end
always @(*) begin
	main_A_a0_a0_in_b = kernel_atax_inst_main_A_a0_a0_in_b;
end
always @(*) begin
	main_A_a0_a0_byteena_b = kernel_atax_inst_main_A_a0_a0_byteena_b;
end
assign main_A_a0_a0_enable_b = 0;
always @(*) begin
	main_A_a0_a0_address_b = kernel_atax_inst_main_A_a0_a0_address_b;
end

endmodule
`timescale 1 ns / 1 ns
module kernel_atax
(
	clk,
	reset,
	start,
	finish,
	main_y_write_enable_a,
	main_y_in_a,
	main_y_byteena_a,
	main_y_enable_a,
	main_y_address_a,
	main_y_out_a,
	main_y_write_enable_b,
	main_y_in_b,
	main_y_byteena_b,
	main_y_enable_b,
	main_y_address_b,
	main_y_out_b,
	main_x_write_enable_a,
	main_x_in_a,
	main_x_byteena_a,
	main_x_enable_a,
	main_x_address_a,
	main_x_out_a,
	main_x_write_enable_b,
	main_x_in_b,
	main_x_byteena_b,
	main_x_enable_b,
	main_x_address_b,
	main_x_out_b,
	main_A_a0_a0_write_enable_a,
	main_A_a0_a0_in_a,
	main_A_a0_a0_byteena_a,
	main_A_a0_a0_enable_a,
	main_A_a0_a0_address_a,
	main_A_a0_a0_out_a,
	main_A_a0_a0_write_enable_b,
	main_A_a0_a0_in_b,
	main_A_a0_a0_byteena_b,
	main_A_a0_a0_enable_b,
	main_A_a0_a0_address_b,
	main_A_a0_a0_out_b
);

parameter [6:0] LEGUP_0 = 7'd0;
parameter [6:0] LEGUP_F_kernel_atax_BB_for_body_1 = 7'd1;
parameter [6:0] LEGUP_F_kernel_atax_BB_for_body_2 = 7'd2;
parameter [6:0] LEGUP_F_kernel_atax_BB_for_body5_preheader_3 = 7'd3;
parameter [6:0] LEGUP_F_kernel_atax_BB_for_body5_4 = 7'd4;
parameter [6:0] LEGUP_F_kernel_atax_BB_for_body9_5 = 7'd5;
parameter [6:0] LEGUP_F_kernel_atax_BB_for_body9_6 = 7'd6;
parameter [6:0] LEGUP_F_kernel_atax_BB_for_body9_7 = 7'd7;
parameter [6:0] LEGUP_F_kernel_atax_BB_for_body9_8 = 7'd8;
parameter [6:0] LEGUP_F_kernel_atax_BB_for_body9_9 = 7'd9;
parameter [6:0] LEGUP_F_kernel_atax_BB_for_body9_10 = 7'd10;
parameter [6:0] LEGUP_F_kernel_atax_BB_for_body9_11 = 7'd11;
parameter [6:0] LEGUP_F_kernel_atax_BB_for_body9_12 = 7'd12;
parameter [6:0] LEGUP_F_kernel_atax_BB_for_body9_13 = 7'd13;
parameter [6:0] LEGUP_F_kernel_atax_BB_for_body9_14 = 7'd14;
parameter [6:0] LEGUP_F_kernel_atax_BB_for_body9_15 = 7'd15;
parameter [6:0] LEGUP_F_kernel_atax_BB_for_body9_16 = 7'd16;
parameter [6:0] LEGUP_F_kernel_atax_BB_for_body9_17 = 7'd17;
parameter [6:0] LEGUP_F_kernel_atax_BB_for_body9_18 = 7'd18;
parameter [6:0] LEGUP_F_kernel_atax_BB_for_body9_19 = 7'd19;
parameter [6:0] LEGUP_F_kernel_atax_BB_for_body9_20 = 7'd20;
parameter [6:0] LEGUP_F_kernel_atax_BB_for_body9_21 = 7'd21;
parameter [6:0] LEGUP_F_kernel_atax_BB_for_body9_22 = 7'd22;
parameter [6:0] LEGUP_F_kernel_atax_BB_for_body9_23 = 7'd23;
parameter [6:0] LEGUP_F_kernel_atax_BB_for_body9_24 = 7'd24;
parameter [6:0] LEGUP_F_kernel_atax_BB_for_body9_25 = 7'd25;
parameter [6:0] LEGUP_F_kernel_atax_BB_for_body9_26 = 7'd26;
parameter [6:0] LEGUP_F_kernel_atax_BB_for_body9_27 = 7'd27;
parameter [6:0] LEGUP_F_kernel_atax_BB_for_body9_28 = 7'd28;
parameter [6:0] LEGUP_F_kernel_atax_BB_for_body9_29 = 7'd29;
parameter [6:0] LEGUP_F_kernel_atax_BB_for_body9_30 = 7'd30;
parameter [6:0] LEGUP_F_kernel_atax_BB_for_body9_31 = 7'd31;
parameter [6:0] LEGUP_F_kernel_atax_BB_for_body9_32 = 7'd32;
parameter [6:0] LEGUP_F_kernel_atax_BB_for_body20_preheader_33 = 7'd33;
parameter [6:0] LEGUP_F_kernel_atax_BB_for_body20_34 = 7'd34;
parameter [6:0] LEGUP_F_kernel_atax_BB_for_body20_35 = 7'd35;
parameter [6:0] LEGUP_F_kernel_atax_BB_for_body20_36 = 7'd36;
parameter [6:0] LEGUP_F_kernel_atax_BB_for_body20_37 = 7'd37;
parameter [6:0] LEGUP_F_kernel_atax_BB_for_body20_38 = 7'd38;
parameter [6:0] LEGUP_F_kernel_atax_BB_for_body20_39 = 7'd39;
parameter [6:0] LEGUP_F_kernel_atax_BB_for_body20_40 = 7'd40;
parameter [6:0] LEGUP_F_kernel_atax_BB_for_body20_41 = 7'd41;
parameter [6:0] LEGUP_F_kernel_atax_BB_for_body20_42 = 7'd42;
parameter [6:0] LEGUP_F_kernel_atax_BB_for_body20_43 = 7'd43;
parameter [6:0] LEGUP_F_kernel_atax_BB_for_body20_44 = 7'd44;
parameter [6:0] LEGUP_F_kernel_atax_BB_for_body20_45 = 7'd45;
parameter [6:0] LEGUP_F_kernel_atax_BB_for_body20_46 = 7'd46;
parameter [6:0] LEGUP_F_kernel_atax_BB_for_body20_47 = 7'd47;
parameter [6:0] LEGUP_F_kernel_atax_BB_for_body20_48 = 7'd48;
parameter [6:0] LEGUP_F_kernel_atax_BB_for_body20_49 = 7'd49;
parameter [6:0] LEGUP_F_kernel_atax_BB_for_body20_50 = 7'd50;
parameter [6:0] LEGUP_F_kernel_atax_BB_for_body20_51 = 7'd51;
parameter [6:0] LEGUP_F_kernel_atax_BB_for_body20_52 = 7'd52;
parameter [6:0] LEGUP_F_kernel_atax_BB_for_body20_53 = 7'd53;
parameter [6:0] LEGUP_F_kernel_atax_BB_for_body20_54 = 7'd54;
parameter [6:0] LEGUP_F_kernel_atax_BB_for_body20_55 = 7'd55;
parameter [6:0] LEGUP_F_kernel_atax_BB_for_body20_56 = 7'd56;
parameter [6:0] LEGUP_F_kernel_atax_BB_for_body20_57 = 7'd57;
parameter [6:0] LEGUP_F_kernel_atax_BB_for_body20_58 = 7'd58;
parameter [6:0] LEGUP_F_kernel_atax_BB_for_body20_59 = 7'd59;
parameter [6:0] LEGUP_F_kernel_atax_BB_for_body20_60 = 7'd60;
parameter [6:0] LEGUP_F_kernel_atax_BB_for_body20_61 = 7'd61;
parameter [6:0] LEGUP_F_kernel_atax_BB_for_body20_62 = 7'd62;
parameter [6:0] LEGUP_F_kernel_atax_BB_for_inc31_63 = 7'd63;
parameter [6:0] LEGUP_F_kernel_atax_BB_for_end33_64 = 7'd64;

input  clk;
input  reset;
input  start;
output reg  finish;
output reg  main_y_write_enable_a;
output reg [63:0] main_y_in_a;
output  main_y_byteena_a;
output reg  main_y_enable_a;
output reg [4:0] main_y_address_a;
input [63:0] main_y_out_a;
output  main_y_write_enable_b;
output [63:0] main_y_in_b;
output  main_y_byteena_b;
output  main_y_enable_b;
output [4:0] main_y_address_b;
input [63:0] main_y_out_b;
output  main_x_write_enable_a;
output [63:0] main_x_in_a;
output  main_x_byteena_a;
output reg  main_x_enable_a;
output reg [4:0] main_x_address_a;
input [63:0] main_x_out_a;
output  main_x_write_enable_b;
output [63:0] main_x_in_b;
output  main_x_byteena_b;
output  main_x_enable_b;
output [4:0] main_x_address_b;
input [63:0] main_x_out_b;
output  main_A_a0_a0_write_enable_a;
output [63:0] main_A_a0_a0_in_a;
output  main_A_a0_a0_byteena_a;
output reg  main_A_a0_a0_enable_a;
output reg [9:0] main_A_a0_a0_address_a;
input [63:0] main_A_a0_a0_out_a;
output  main_A_a0_a0_write_enable_b;
output [63:0] main_A_a0_a0_in_b;
output  main_A_a0_a0_byteena_b;
output  main_A_a0_a0_enable_b;
output [9:0] main_A_a0_a0_address_b;
input [63:0] main_A_a0_a0_out_b;
reg [6:0] cur_state;
reg [6:0] next_state;
wire  fsm_stall;
reg [5:0] kernel_atax_for_body_i_04;
reg [5:0] kernel_atax_for_body_i_04_reg;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] kernel_atax_for_body_arrayidx;
reg [6:0] kernel_atax_for_body_0;
reg [6:0] kernel_atax_for_body_0_reg;
reg  kernel_atax_for_body_exitcond13;
reg  kernel_atax_for_body_exitcond13_reg;
reg [5:0] kernel_atax_for_body5_i_13;
reg [5:0] kernel_atax_for_body5_i_13_reg;
reg [26:0] kernel_atax_for_body5_bit_select;
reg [31:0] kernel_atax_for_body5_bit_concat;
reg [31:0] kernel_atax_for_body5_bit_concat_reg;
reg [63:0] kernel_atax_for_body9_1;
reg [63:0] kernel_atax_for_body9_1_reg;
reg [31:0] kernel_atax_for_body9_j_01;
reg [31:0] kernel_atax_for_body9_j_01_reg;
reg [31:0] kernel_atax_for_body9_2;
reg [31:0] kernel_atax_for_body9_2_reg;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] kernel_atax_for_body9_scevgep;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] kernel_atax_for_body9_arrayidx13;
reg [63:0] kernel_atax_for_body9_3;
reg [63:0] kernel_atax_for_body9_4;
reg [63:0] kernel_atax_for_body9_4_reg;
reg [63:0] kernel_atax_for_body9_mul;
reg [63:0] kernel_atax_for_body9_add;
reg [63:0] kernel_atax_for_body9_add_reg;
reg [31:0] kernel_atax_for_body9_5;
reg [31:0] kernel_atax_for_body9_5_reg;
reg  kernel_atax_for_body9_exitcond3;
reg  kernel_atax_for_body9_exitcond3_reg;
reg [31:0] kernel_atax_for_body20_j_12;
reg [31:0] kernel_atax_for_body20_j_12_reg;
reg [31:0] kernel_atax_for_body20_6;
reg [31:0] kernel_atax_for_body20_6_reg;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] kernel_atax_for_body20_scevgep4;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] kernel_atax_for_body20_arrayidx21;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] kernel_atax_for_body20_arrayidx21_reg;
reg [63:0] kernel_atax_for_body20_7;
reg [63:0] kernel_atax_for_body20_7_reg;
reg [63:0] kernel_atax_for_body20_8;
reg [63:0] kernel_atax_for_body20_mul25;
reg [63:0] kernel_atax_for_body20_add26;
reg [31:0] kernel_atax_for_body20_9;
reg [31:0] kernel_atax_for_body20_9_reg;
reg  kernel_atax_for_body20_exitcond7;
reg  kernel_atax_for_body20_exitcond7_reg;
reg [6:0] kernel_atax_for_inc31_10;
reg  kernel_atax_for_inc31_exitcond10;
reg [63:0] kernel_atax_altfp_multiply_64_0_op0;
reg [63:0] kernel_atax_altfp_multiply_64_0_op1;
reg  kernel_atax_altfp_multiply_64_0_inst_clock;
reg  kernel_atax_altfp_multiply_64_0_inst_clk_en;
reg [63:0] kernel_atax_altfp_multiply_64_0_inst_dataa;
reg [63:0] kernel_atax_altfp_multiply_64_0_inst_datab;
wire [63:0] kernel_atax_altfp_multiply_64_0_inst_result;
reg [63:0] kernel_atax_for_body9_mul_out;
reg  altfp_kernel_atax_for_body9_mul_en;
reg [63:0] kernel_atax_altfp_multiply_64_0;
reg [63:0] kernel_atax_altfp_add_64_0_op0;
reg [63:0] kernel_atax_altfp_add_64_0_op1;
reg  kernel_atax_altfp_add_64_0_inst_clock;
reg  kernel_atax_altfp_add_64_0_inst_clk_en;
reg [63:0] kernel_atax_altfp_add_64_0_inst_dataa;
reg [63:0] kernel_atax_altfp_add_64_0_inst_datab;
wire [63:0] kernel_atax_altfp_add_64_0_inst_result;
reg [63:0] kernel_atax_for_body9_add_out;
reg  altfp_kernel_atax_for_body9_add_en;
reg [63:0] kernel_atax_altfp_add_64_0;
reg [26:0] kernel_atax_for_body5_i_13_reg_width_extended;
wire [4:0] kernel_atax_for_body5_bit_concat_bit_select_operand_2;


altfp_multiplier64_11 kernel_atax_altfp_multiply_64_0_inst (
	.clock (kernel_atax_altfp_multiply_64_0_inst_clock),
	.clk_en (kernel_atax_altfp_multiply_64_0_inst_clk_en),
	.dataa (kernel_atax_altfp_multiply_64_0_inst_dataa),
	.datab (kernel_atax_altfp_multiply_64_0_inst_datab),
	.result (kernel_atax_altfp_multiply_64_0_inst_result)
);



altfp_adder64_14 kernel_atax_altfp_add_64_0_inst (
	.clock (kernel_atax_altfp_add_64_0_inst_clock),
	.clk_en (kernel_atax_altfp_add_64_0_inst_clk_en),
	.dataa (kernel_atax_altfp_add_64_0_inst_dataa),
	.datab (kernel_atax_altfp_add_64_0_inst_datab),
	.result (kernel_atax_altfp_add_64_0_inst_result)
);



always @(posedge clk) begin
if (reset == 1'b1)
	cur_state <= LEGUP_0;
else if (!fsm_stall)
	cur_state <= next_state;
end

always @(*)
begin
next_state = cur_state;
case(cur_state)  // synthesis parallel_case  
LEGUP_0:
	if ((fsm_stall == 1'd0) && (start == 1'd1))
		next_state = LEGUP_F_kernel_atax_BB_for_body_1;
LEGUP_F_kernel_atax_BB_for_body20_34:
		next_state = LEGUP_F_kernel_atax_BB_for_body20_35;
LEGUP_F_kernel_atax_BB_for_body20_35:
		next_state = LEGUP_F_kernel_atax_BB_for_body20_36;
LEGUP_F_kernel_atax_BB_for_body20_36:
		next_state = LEGUP_F_kernel_atax_BB_for_body20_37;
LEGUP_F_kernel_atax_BB_for_body20_37:
		next_state = LEGUP_F_kernel_atax_BB_for_body20_38;
LEGUP_F_kernel_atax_BB_for_body20_38:
		next_state = LEGUP_F_kernel_atax_BB_for_body20_39;
LEGUP_F_kernel_atax_BB_for_body20_39:
		next_state = LEGUP_F_kernel_atax_BB_for_body20_40;
LEGUP_F_kernel_atax_BB_for_body20_40:
		next_state = LEGUP_F_kernel_atax_BB_for_body20_41;
LEGUP_F_kernel_atax_BB_for_body20_41:
		next_state = LEGUP_F_kernel_atax_BB_for_body20_42;
LEGUP_F_kernel_atax_BB_for_body20_42:
		next_state = LEGUP_F_kernel_atax_BB_for_body20_43;
LEGUP_F_kernel_atax_BB_for_body20_43:
		next_state = LEGUP_F_kernel_atax_BB_for_body20_44;
LEGUP_F_kernel_atax_BB_for_body20_44:
		next_state = LEGUP_F_kernel_atax_BB_for_body20_45;
LEGUP_F_kernel_atax_BB_for_body20_45:
		next_state = LEGUP_F_kernel_atax_BB_for_body20_46;
LEGUP_F_kernel_atax_BB_for_body20_46:
		next_state = LEGUP_F_kernel_atax_BB_for_body20_47;
LEGUP_F_kernel_atax_BB_for_body20_47:
		next_state = LEGUP_F_kernel_atax_BB_for_body20_48;
LEGUP_F_kernel_atax_BB_for_body20_48:
		next_state = LEGUP_F_kernel_atax_BB_for_body20_49;
LEGUP_F_kernel_atax_BB_for_body20_49:
		next_state = LEGUP_F_kernel_atax_BB_for_body20_50;
LEGUP_F_kernel_atax_BB_for_body20_50:
		next_state = LEGUP_F_kernel_atax_BB_for_body20_51;
LEGUP_F_kernel_atax_BB_for_body20_51:
		next_state = LEGUP_F_kernel_atax_BB_for_body20_52;
LEGUP_F_kernel_atax_BB_for_body20_52:
		next_state = LEGUP_F_kernel_atax_BB_for_body20_53;
LEGUP_F_kernel_atax_BB_for_body20_53:
		next_state = LEGUP_F_kernel_atax_BB_for_body20_54;
LEGUP_F_kernel_atax_BB_for_body20_54:
		next_state = LEGUP_F_kernel_atax_BB_for_body20_55;
LEGUP_F_kernel_atax_BB_for_body20_55:
		next_state = LEGUP_F_kernel_atax_BB_for_body20_56;
LEGUP_F_kernel_atax_BB_for_body20_56:
		next_state = LEGUP_F_kernel_atax_BB_for_body20_57;
LEGUP_F_kernel_atax_BB_for_body20_57:
		next_state = LEGUP_F_kernel_atax_BB_for_body20_58;
LEGUP_F_kernel_atax_BB_for_body20_58:
		next_state = LEGUP_F_kernel_atax_BB_for_body20_59;
LEGUP_F_kernel_atax_BB_for_body20_59:
		next_state = LEGUP_F_kernel_atax_BB_for_body20_60;
LEGUP_F_kernel_atax_BB_for_body20_60:
		next_state = LEGUP_F_kernel_atax_BB_for_body20_61;
LEGUP_F_kernel_atax_BB_for_body20_61:
		next_state = LEGUP_F_kernel_atax_BB_for_body20_62;
LEGUP_F_kernel_atax_BB_for_body20_62:
	if ((fsm_stall == 1'd0) && (kernel_atax_for_body20_exitcond7_reg == 1'd1))
		next_state = LEGUP_F_kernel_atax_BB_for_inc31_63;
	else if ((fsm_stall == 1'd0) && (kernel_atax_for_body20_exitcond7_reg == 1'd0))
		next_state = LEGUP_F_kernel_atax_BB_for_body20_34;
LEGUP_F_kernel_atax_BB_for_body20_preheader_33:
		next_state = LEGUP_F_kernel_atax_BB_for_body20_34;
LEGUP_F_kernel_atax_BB_for_body5_4:
		next_state = LEGUP_F_kernel_atax_BB_for_body9_5;
LEGUP_F_kernel_atax_BB_for_body5_preheader_3:
		next_state = LEGUP_F_kernel_atax_BB_for_body5_4;
LEGUP_F_kernel_atax_BB_for_body9_10:
		next_state = LEGUP_F_kernel_atax_BB_for_body9_11;
LEGUP_F_kernel_atax_BB_for_body9_11:
		next_state = LEGUP_F_kernel_atax_BB_for_body9_12;
LEGUP_F_kernel_atax_BB_for_body9_12:
		next_state = LEGUP_F_kernel_atax_BB_for_body9_13;
LEGUP_F_kernel_atax_BB_for_body9_13:
		next_state = LEGUP_F_kernel_atax_BB_for_body9_14;
LEGUP_F_kernel_atax_BB_for_body9_14:
		next_state = LEGUP_F_kernel_atax_BB_for_body9_15;
LEGUP_F_kernel_atax_BB_for_body9_15:
		next_state = LEGUP_F_kernel_atax_BB_for_body9_16;
LEGUP_F_kernel_atax_BB_for_body9_16:
		next_state = LEGUP_F_kernel_atax_BB_for_body9_17;
LEGUP_F_kernel_atax_BB_for_body9_17:
		next_state = LEGUP_F_kernel_atax_BB_for_body9_18;
LEGUP_F_kernel_atax_BB_for_body9_18:
		next_state = LEGUP_F_kernel_atax_BB_for_body9_19;
LEGUP_F_kernel_atax_BB_for_body9_19:
		next_state = LEGUP_F_kernel_atax_BB_for_body9_20;
LEGUP_F_kernel_atax_BB_for_body9_20:
		next_state = LEGUP_F_kernel_atax_BB_for_body9_21;
LEGUP_F_kernel_atax_BB_for_body9_21:
		next_state = LEGUP_F_kernel_atax_BB_for_body9_22;
LEGUP_F_kernel_atax_BB_for_body9_22:
		next_state = LEGUP_F_kernel_atax_BB_for_body9_23;
LEGUP_F_kernel_atax_BB_for_body9_23:
		next_state = LEGUP_F_kernel_atax_BB_for_body9_24;
LEGUP_F_kernel_atax_BB_for_body9_24:
		next_state = LEGUP_F_kernel_atax_BB_for_body9_25;
LEGUP_F_kernel_atax_BB_for_body9_25:
		next_state = LEGUP_F_kernel_atax_BB_for_body9_26;
LEGUP_F_kernel_atax_BB_for_body9_26:
		next_state = LEGUP_F_kernel_atax_BB_for_body9_27;
LEGUP_F_kernel_atax_BB_for_body9_27:
		next_state = LEGUP_F_kernel_atax_BB_for_body9_28;
LEGUP_F_kernel_atax_BB_for_body9_28:
		next_state = LEGUP_F_kernel_atax_BB_for_body9_29;
LEGUP_F_kernel_atax_BB_for_body9_29:
		next_state = LEGUP_F_kernel_atax_BB_for_body9_30;
LEGUP_F_kernel_atax_BB_for_body9_30:
		next_state = LEGUP_F_kernel_atax_BB_for_body9_31;
LEGUP_F_kernel_atax_BB_for_body9_31:
		next_state = LEGUP_F_kernel_atax_BB_for_body9_32;
LEGUP_F_kernel_atax_BB_for_body9_32:
	if ((fsm_stall == 1'd0) && (kernel_atax_for_body9_exitcond3_reg == 1'd1))
		next_state = LEGUP_F_kernel_atax_BB_for_body20_preheader_33;
	else if ((fsm_stall == 1'd0) && (kernel_atax_for_body9_exitcond3_reg == 1'd0))
		next_state = LEGUP_F_kernel_atax_BB_for_body9_5;
LEGUP_F_kernel_atax_BB_for_body9_5:
		next_state = LEGUP_F_kernel_atax_BB_for_body9_6;
LEGUP_F_kernel_atax_BB_for_body9_6:
		next_state = LEGUP_F_kernel_atax_BB_for_body9_7;
LEGUP_F_kernel_atax_BB_for_body9_7:
		next_state = LEGUP_F_kernel_atax_BB_for_body9_8;
LEGUP_F_kernel_atax_BB_for_body9_8:
		next_state = LEGUP_F_kernel_atax_BB_for_body9_9;
LEGUP_F_kernel_atax_BB_for_body9_9:
		next_state = LEGUP_F_kernel_atax_BB_for_body9_10;
LEGUP_F_kernel_atax_BB_for_body_1:
		next_state = LEGUP_F_kernel_atax_BB_for_body_2;
LEGUP_F_kernel_atax_BB_for_body_2:
	if ((fsm_stall == 1'd0) && (kernel_atax_for_body_exitcond13_reg == 1'd1))
		next_state = LEGUP_F_kernel_atax_BB_for_body5_preheader_3;
	else if ((fsm_stall == 1'd0) && (kernel_atax_for_body_exitcond13_reg == 1'd0))
		next_state = LEGUP_F_kernel_atax_BB_for_body_1;
LEGUP_F_kernel_atax_BB_for_end33_64:
		next_state = LEGUP_0;
LEGUP_F_kernel_atax_BB_for_inc31_63:
	if ((fsm_stall == 1'd0) && (kernel_atax_for_inc31_exitcond10 == 1'd1))
		next_state = LEGUP_F_kernel_atax_BB_for_end33_64;
	else if ((fsm_stall == 1'd0) && (kernel_atax_for_inc31_exitcond10 == 1'd0))
		next_state = LEGUP_F_kernel_atax_BB_for_body5_4;
default:
	next_state = cur_state;
endcase

end
assign fsm_stall = 1'd0;
always @(*) begin
	if ((((cur_state == LEGUP_0) & (fsm_stall == 1'd0)) & (start == 1'd1))) begin
		kernel_atax_for_body_i_04 = 32'd0;
	end
	else /* if ((((cur_state == LEGUP_F_kernel_atax_BB_for_body_2) & (fsm_stall == 1'd0)) & (kernel_atax_for_body_exitcond13_reg == 1'd0))) */ begin
		kernel_atax_for_body_i_04 = kernel_atax_for_body_0_reg;
	end
end
always @(posedge clk) begin
	if ((((cur_state == LEGUP_0) & (fsm_stall == 1'd0)) & (start == 1'd1))) begin
		kernel_atax_for_body_i_04_reg <= kernel_atax_for_body_i_04;
	end
	if ((((cur_state == LEGUP_F_kernel_atax_BB_for_body_2) & (fsm_stall == 1'd0)) & (kernel_atax_for_body_exitcond13_reg == 1'd0))) begin
		kernel_atax_for_body_i_04_reg <= kernel_atax_for_body_i_04;
	end
end
always @(*) begin
		kernel_atax_for_body_arrayidx = (1'd0 + (8 * {26'd0,kernel_atax_for_body_i_04_reg}));
end
always @(*) begin
		kernel_atax_for_body_0 = ({1'd0,kernel_atax_for_body_i_04_reg} + 32'd1);
end
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_kernel_atax_BB_for_body_1)) begin
		kernel_atax_for_body_0_reg <= kernel_atax_for_body_0;
	end
end
always @(*) begin
		kernel_atax_for_body_exitcond13 = (kernel_atax_for_body_0 == 32'd32);
end
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_kernel_atax_BB_for_body_1)) begin
		kernel_atax_for_body_exitcond13_reg <= kernel_atax_for_body_exitcond13;
	end
end
always @(*) begin
	if (((cur_state == LEGUP_F_kernel_atax_BB_for_body5_preheader_3) & (fsm_stall == 1'd0))) begin
		kernel_atax_for_body5_i_13 = 32'd0;
	end
	else /* if ((((cur_state == LEGUP_F_kernel_atax_BB_for_inc31_63) & (fsm_stall == 1'd0)) & (kernel_atax_for_inc31_exitcond10 == 1'd0))) */ begin
		kernel_atax_for_body5_i_13 = kernel_atax_for_inc31_10;
	end
end
always @(posedge clk) begin
	if (((cur_state == LEGUP_F_kernel_atax_BB_for_body5_preheader_3) & (fsm_stall == 1'd0))) begin
		kernel_atax_for_body5_i_13_reg <= kernel_atax_for_body5_i_13;
	end
	if ((((cur_state == LEGUP_F_kernel_atax_BB_for_inc31_63) & (fsm_stall == 1'd0)) & (kernel_atax_for_inc31_exitcond10 == 1'd0))) begin
		kernel_atax_for_body5_i_13_reg <= kernel_atax_for_body5_i_13;
	end
end
always @(*) begin
		kernel_atax_for_body5_bit_select = kernel_atax_for_body5_i_13_reg_width_extended[26:0];
end
always @(*) begin
		kernel_atax_for_body5_bit_concat = {kernel_atax_for_body5_bit_select[26:0], kernel_atax_for_body5_bit_concat_bit_select_operand_2[4:0]};
end
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_kernel_atax_BB_for_body5_4)) begin
		kernel_atax_for_body5_bit_concat_reg <= kernel_atax_for_body5_bit_concat;
	end
end
always @(*) begin
	if (((cur_state == LEGUP_F_kernel_atax_BB_for_body5_4) & (fsm_stall == 1'd0))) begin
		kernel_atax_for_body9_1 = 64'h0;
	end
	else /* if ((((cur_state == LEGUP_F_kernel_atax_BB_for_body9_32) & (fsm_stall == 1'd0)) & (kernel_atax_for_body9_exitcond3_reg == 1'd0))) */ begin
		kernel_atax_for_body9_1 = kernel_atax_for_body9_add;
	end
end
always @(posedge clk) begin
	if (((cur_state == LEGUP_F_kernel_atax_BB_for_body5_4) & (fsm_stall == 1'd0))) begin
		kernel_atax_for_body9_1_reg <= kernel_atax_for_body9_1;
	end
	if ((((cur_state == LEGUP_F_kernel_atax_BB_for_body9_32) & (fsm_stall == 1'd0)) & (kernel_atax_for_body9_exitcond3_reg == 1'd0))) begin
		kernel_atax_for_body9_1_reg <= kernel_atax_for_body9_1;
	end
end
always @(*) begin
	if (((cur_state == LEGUP_F_kernel_atax_BB_for_body5_4) & (fsm_stall == 1'd0))) begin
		kernel_atax_for_body9_j_01 = 32'd0;
	end
	else /* if ((((cur_state == LEGUP_F_kernel_atax_BB_for_body9_32) & (fsm_stall == 1'd0)) & (kernel_atax_for_body9_exitcond3_reg == 1'd0))) */ begin
		kernel_atax_for_body9_j_01 = kernel_atax_for_body9_5_reg;
	end
end
always @(posedge clk) begin
	if (((cur_state == LEGUP_F_kernel_atax_BB_for_body5_4) & (fsm_stall == 1'd0))) begin
		kernel_atax_for_body9_j_01_reg <= kernel_atax_for_body9_j_01;
	end
	if ((((cur_state == LEGUP_F_kernel_atax_BB_for_body9_32) & (fsm_stall == 1'd0)) & (kernel_atax_for_body9_exitcond3_reg == 1'd0))) begin
		kernel_atax_for_body9_j_01_reg <= kernel_atax_for_body9_j_01;
	end
end
always @(*) begin
		kernel_atax_for_body9_2 = (kernel_atax_for_body5_bit_concat_reg + kernel_atax_for_body9_j_01_reg);
end
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_kernel_atax_BB_for_body9_5)) begin
		kernel_atax_for_body9_2_reg <= kernel_atax_for_body9_2;
	end
end
always @(*) begin
		kernel_atax_for_body9_scevgep = (1'd0 + (8 * kernel_atax_for_body9_2_reg));
end
always @(*) begin
		kernel_atax_for_body9_arrayidx13 = (1'd0 + (8 * kernel_atax_for_body9_j_01_reg));
end
always @(*) begin
		kernel_atax_for_body9_3 = main_A_a0_a0_out_a;
end
always @(*) begin
		kernel_atax_for_body9_4 = main_x_out_a;
end
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_kernel_atax_BB_for_body9_6)) begin
		kernel_atax_for_body9_4_reg <= kernel_atax_for_body9_4;
	end
end
always @(*) begin
	kernel_atax_for_body9_mul = kernel_atax_altfp_multiply_64_0;
end
always @(*) begin
	kernel_atax_for_body9_add = kernel_atax_altfp_add_64_0;
end
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_kernel_atax_BB_for_body9_32)) begin
		kernel_atax_for_body9_add_reg <= kernel_atax_for_body9_add;
	end
end
always @(*) begin
		kernel_atax_for_body9_5 = (kernel_atax_for_body9_j_01_reg + 32'd1);
end
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_kernel_atax_BB_for_body9_5)) begin
		kernel_atax_for_body9_5_reg <= kernel_atax_for_body9_5;
	end
end
always @(*) begin
		kernel_atax_for_body9_exitcond3 = (kernel_atax_for_body9_5 == 32'd32);
end
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_kernel_atax_BB_for_body9_5)) begin
		kernel_atax_for_body9_exitcond3_reg <= kernel_atax_for_body9_exitcond3;
	end
end
always @(*) begin
	if (((cur_state == LEGUP_F_kernel_atax_BB_for_body20_preheader_33) & (fsm_stall == 1'd0))) begin
		kernel_atax_for_body20_j_12 = 32'd0;
	end
	else /* if ((((cur_state == LEGUP_F_kernel_atax_BB_for_body20_62) & (fsm_stall == 1'd0)) & (kernel_atax_for_body20_exitcond7_reg == 1'd0))) */ begin
		kernel_atax_for_body20_j_12 = kernel_atax_for_body20_9_reg;
	end
end
always @(posedge clk) begin
	if (((cur_state == LEGUP_F_kernel_atax_BB_for_body20_preheader_33) & (fsm_stall == 1'd0))) begin
		kernel_atax_for_body20_j_12_reg <= kernel_atax_for_body20_j_12;
	end
	if ((((cur_state == LEGUP_F_kernel_atax_BB_for_body20_62) & (fsm_stall == 1'd0)) & (kernel_atax_for_body20_exitcond7_reg == 1'd0))) begin
		kernel_atax_for_body20_j_12_reg <= kernel_atax_for_body20_j_12;
	end
end
always @(*) begin
		kernel_atax_for_body20_6 = (kernel_atax_for_body5_bit_concat_reg + kernel_atax_for_body20_j_12_reg);
end
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_kernel_atax_BB_for_body20_34)) begin
		kernel_atax_for_body20_6_reg <= kernel_atax_for_body20_6;
	end
end
always @(*) begin
		kernel_atax_for_body20_scevgep4 = (1'd0 + (8 * kernel_atax_for_body20_6_reg));
end
always @(*) begin
		kernel_atax_for_body20_arrayidx21 = (1'd0 + (8 * kernel_atax_for_body20_j_12_reg));
end
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_kernel_atax_BB_for_body20_34)) begin
		kernel_atax_for_body20_arrayidx21_reg <= kernel_atax_for_body20_arrayidx21;
	end
end
always @(*) begin
		kernel_atax_for_body20_7 = main_y_out_a;
end
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_kernel_atax_BB_for_body20_35)) begin
		kernel_atax_for_body20_7_reg <= kernel_atax_for_body20_7;
	end
end
always @(*) begin
		kernel_atax_for_body20_8 = main_A_a0_a0_out_a;
end
always @(*) begin
	kernel_atax_for_body20_mul25 = kernel_atax_altfp_multiply_64_0;
end
always @(*) begin
	kernel_atax_for_body20_add26 = kernel_atax_altfp_add_64_0;
end
always @(*) begin
		kernel_atax_for_body20_9 = (kernel_atax_for_body20_j_12_reg + 32'd1);
end
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_kernel_atax_BB_for_body20_34)) begin
		kernel_atax_for_body20_9_reg <= kernel_atax_for_body20_9;
	end
end
always @(*) begin
		kernel_atax_for_body20_exitcond7 = (kernel_atax_for_body20_9 == 32'd32);
end
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_kernel_atax_BB_for_body20_34)) begin
		kernel_atax_for_body20_exitcond7_reg <= kernel_atax_for_body20_exitcond7;
	end
end
always @(*) begin
		kernel_atax_for_inc31_10 = ({1'd0,kernel_atax_for_body5_i_13_reg} + 32'd1);
end
always @(*) begin
		kernel_atax_for_inc31_exitcond10 = (kernel_atax_for_inc31_10 == 32'd32);
end
always @(*) begin
	if ((cur_state == LEGUP_F_kernel_atax_BB_for_body9_7)) begin
		kernel_atax_altfp_multiply_64_0_op0 = kernel_atax_for_body9_3;
	end
	else /* if ((cur_state == LEGUP_F_kernel_atax_BB_for_body20_36)) */ begin
		kernel_atax_altfp_multiply_64_0_op0 = kernel_atax_for_body20_8;
	end
end
always @(*) begin
	if ((cur_state == LEGUP_F_kernel_atax_BB_for_body9_7)) begin
		kernel_atax_altfp_multiply_64_0_op1 = kernel_atax_for_body9_4_reg;
	end
	else /* if ((cur_state == LEGUP_F_kernel_atax_BB_for_body20_36)) */ begin
		kernel_atax_altfp_multiply_64_0_op1 = kernel_atax_for_body9_add_reg;
	end
end
always @(*) begin
	kernel_atax_altfp_multiply_64_0_inst_clock = clk;
end
always @(*) begin
	kernel_atax_altfp_multiply_64_0_inst_clk_en = altfp_kernel_atax_for_body9_mul_en;
end
always @(*) begin
	kernel_atax_altfp_multiply_64_0_inst_dataa = kernel_atax_altfp_multiply_64_0_op0;
end
always @(*) begin
	kernel_atax_altfp_multiply_64_0_inst_datab = kernel_atax_altfp_multiply_64_0_op1;
end
always @(*) begin
	kernel_atax_for_body9_mul_out = kernel_atax_altfp_multiply_64_0_inst_result;
end
always @(*) begin
	altfp_kernel_atax_for_body9_mul_en = ~(fsm_stall);
end
always @(*) begin
	kernel_atax_altfp_multiply_64_0 = kernel_atax_for_body9_mul_out;
end
always @(*) begin
	if ((cur_state == LEGUP_F_kernel_atax_BB_for_body9_18)) begin
		kernel_atax_altfp_add_64_0_op0 = kernel_atax_for_body9_1_reg;
	end
	else /* if ((cur_state == LEGUP_F_kernel_atax_BB_for_body20_47)) */ begin
		kernel_atax_altfp_add_64_0_op0 = kernel_atax_for_body20_7_reg;
	end
end
always @(*) begin
	if ((cur_state == LEGUP_F_kernel_atax_BB_for_body9_18)) begin
		kernel_atax_altfp_add_64_0_op1 = kernel_atax_for_body9_mul;
	end
	else /* if ((cur_state == LEGUP_F_kernel_atax_BB_for_body20_47)) */ begin
		kernel_atax_altfp_add_64_0_op1 = kernel_atax_for_body20_mul25;
	end
end
always @(*) begin
	kernel_atax_altfp_add_64_0_inst_clock = clk;
end
always @(*) begin
	kernel_atax_altfp_add_64_0_inst_clk_en = altfp_kernel_atax_for_body9_add_en;
end
always @(*) begin
	kernel_atax_altfp_add_64_0_inst_dataa = kernel_atax_altfp_add_64_0_op0;
end
always @(*) begin
	kernel_atax_altfp_add_64_0_inst_datab = kernel_atax_altfp_add_64_0_op1;
end
always @(*) begin
	kernel_atax_for_body9_add_out = kernel_atax_altfp_add_64_0_inst_result;
end
always @(*) begin
	altfp_kernel_atax_for_body9_add_en = ~(fsm_stall);
end
always @(*) begin
	kernel_atax_altfp_add_64_0 = kernel_atax_for_body9_add_out;
end
always @(*) begin
	kernel_atax_for_body5_i_13_reg_width_extended = {21'd0,kernel_atax_for_body5_i_13_reg};
end
assign kernel_atax_for_body5_bit_concat_bit_select_operand_2 = 5'd0;
always @(posedge clk) begin
	if ((cur_state == LEGUP_0)) begin
		finish <= 1'd0;
	end
	if ((cur_state == LEGUP_F_kernel_atax_BB_for_end33_64)) begin
		finish <= (fsm_stall == 1'd0);
	end
end
always @(*) begin
	main_y_write_enable_a = 1'd0;
	if ((cur_state == LEGUP_F_kernel_atax_BB_for_body_1)) begin
		main_y_write_enable_a = 1'd1;
	end
	if ((cur_state == LEGUP_F_kernel_atax_BB_for_body20_61)) begin
		main_y_write_enable_a = 1'd1;
	end
end
always @(*) begin
	main_y_in_a = 64'd0;
	if ((cur_state == LEGUP_F_kernel_atax_BB_for_body_1)) begin
		main_y_in_a = 64'h0;
	end
	if ((cur_state == LEGUP_F_kernel_atax_BB_for_body20_61)) begin
		main_y_in_a = kernel_atax_for_body20_add26;
	end
end
assign main_y_byteena_a = 1'd1;
always @(*) begin
	main_y_enable_a = 1'd0;
	if ((cur_state == LEGUP_F_kernel_atax_BB_for_body_1)) begin
		main_y_enable_a = 1'd1;
	end
	if ((cur_state == LEGUP_F_kernel_atax_BB_for_body20_34)) begin
		main_y_enable_a = 1'd1;
	end
	if ((cur_state == LEGUP_F_kernel_atax_BB_for_body20_61)) begin
		main_y_enable_a = 1'd1;
	end
end
always @(*) begin
	main_y_address_a = 5'd0;
	if ((cur_state == LEGUP_F_kernel_atax_BB_for_body_1)) begin
		main_y_address_a = (kernel_atax_for_body_arrayidx >>> 3'd3);
	end
	if ((cur_state == LEGUP_F_kernel_atax_BB_for_body20_34)) begin
		main_y_address_a = (kernel_atax_for_body20_arrayidx21 >>> 3'd3);
	end
	if ((cur_state == LEGUP_F_kernel_atax_BB_for_body20_61)) begin
		main_y_address_a = (kernel_atax_for_body20_arrayidx21_reg >>> 3'd3);
	end
end
assign main_y_write_enable_b = 1'd0;
assign main_y_in_b = 64'd0;
assign main_y_byteena_b = 1'd1;
assign main_y_enable_b = 1'd0;
assign main_y_address_b = 5'd0;
assign main_x_write_enable_a = 1'd0;
assign main_x_in_a = 64'd0;
assign main_x_byteena_a = 1'd1;
always @(*) begin
	main_x_enable_a = 1'd0;
	if ((cur_state == LEGUP_F_kernel_atax_BB_for_body9_5)) begin
		main_x_enable_a = 1'd1;
	end
end
always @(*) begin
	main_x_address_a = 5'd0;
	if ((cur_state == LEGUP_F_kernel_atax_BB_for_body9_5)) begin
		main_x_address_a = (kernel_atax_for_body9_arrayidx13 >>> 3'd3);
	end
end
assign main_x_write_enable_b = 1'd0;
assign main_x_in_b = 64'd0;
assign main_x_byteena_b = 1'd1;
assign main_x_enable_b = 1'd0;
assign main_x_address_b = 5'd0;
assign main_A_a0_a0_write_enable_a = 1'd0;
assign main_A_a0_a0_in_a = 64'd0;
assign main_A_a0_a0_byteena_a = 1'd1;
always @(*) begin
	main_A_a0_a0_enable_a = 1'd0;
	if ((cur_state == LEGUP_F_kernel_atax_BB_for_body9_6)) begin
		main_A_a0_a0_enable_a = 1'd1;
	end
	if ((cur_state == LEGUP_F_kernel_atax_BB_for_body20_35)) begin
		main_A_a0_a0_enable_a = 1'd1;
	end
end
always @(*) begin
	main_A_a0_a0_address_a = 10'd0;
	if ((cur_state == LEGUP_F_kernel_atax_BB_for_body9_6)) begin
		main_A_a0_a0_address_a = (kernel_atax_for_body9_scevgep >>> 3'd3);
	end
	if ((cur_state == LEGUP_F_kernel_atax_BB_for_body20_35)) begin
		main_A_a0_a0_address_a = (kernel_atax_for_body20_scevgep4 >>> 3'd3);
	end
end
assign main_A_a0_a0_write_enable_b = 1'd0;
assign main_A_a0_a0_in_b = 64'd0;
assign main_A_a0_a0_byteena_b = 1'd1;
assign main_A_a0_a0_enable_b = 1'd0;
assign main_A_a0_a0_address_b = 10'd0;

endmodule


module ram_dual_port
(
	clk,
	clken,
	address_a,
	address_b,
	wren_a,
	data_a,
	byteena_a,
	wren_b,
	data_b,
	byteena_b,
	q_b,
	q_a
);

parameter  width_a = 1'd0;
parameter  widthad_a = 1'd0;
parameter  numwords_a = 1'd0;
parameter  width_b = 1'd0;
parameter  widthad_b = 1'd0;
parameter  numwords_b = 1'd0;
parameter  latency = 1;
parameter  init_file = "UNUSED";
parameter  width_be_a = 1'd0;
parameter  width_be_b = 1'd0;
localparam output_registered = (latency == 1)? "UNREGISTERED" : "CLOCK0";
input  clk;
input  clken;
input [(widthad_a-1):0] address_a;
output wire [(width_a-1):0] q_a;
wire [(width_a-1):0] q_a_wire;
input [(widthad_b-1):0] address_b;
output wire [(width_b-1):0] q_b;
wire [(width_b-1):0] q_b_wire;
input  wren_a;
input [(width_a-1):0] data_a;
input [width_be_a-1:0] byteena_a;
input  wren_b;
input [(width_b-1):0] data_b;
input [width_be_b-1:0] byteena_b;
reg  clk_wire;

altsyncram altsyncram_component (
	.address_a (address_a),
    .clock0 (clk_wire),
    .clock1 (1'd1),
    .clocken0 (clken),
    .clocken1 (1'd1),
    .clocken2 (1'd1),
    .clocken3 (1'd1),
    .aclr0 (1'd0),
    .aclr1 (1'd0),
    .addressstall_a (1'd0),
    .eccstatus (),
    .rden_a (clken),
    .q_a (q_a),
	.address_b (address_b),
    .addressstall_b (1'd0),
    .rden_b (clken),
    .q_b (q_b),
    .wren_a (wren_a),
    .data_a (data_a),
    .wren_b (wren_b),
    .data_b (data_b),
    .byteena_b (byteena_b),
    .byteena_a (byteena_a)
);
defparam
    altsyncram_component.width_byteena_a = width_be_a,
    altsyncram_component.width_byteena_b = width_be_b,
    altsyncram_component.operation_mode = "BIDIR_DUAL_PORT",
    altsyncram_component.read_during_write_mode_mixed_ports = "OLD_DATA",
    altsyncram_component.init_file = init_file,
    altsyncram_component.lpm_hint = "ENABLE_RUNTIME_MOD=NO",
    altsyncram_component.lpm_type = "altsyncram",
    altsyncram_component.power_up_uninitialized = "FALSE",
    altsyncram_component.intended_device_family = "CycloneV",
    altsyncram_component.clock_enable_input_b = "BYPASS",
    altsyncram_component.clock_enable_output_b = "BYPASS",
    altsyncram_component.outdata_aclr_b = "NONE",
    altsyncram_component.outdata_reg_b = output_registered,
    altsyncram_component.numwords_b = numwords_b,
    altsyncram_component.widthad_b = widthad_b,
    altsyncram_component.width_b = width_b,
    altsyncram_component.address_reg_b = "CLOCK0",
    altsyncram_component.byteena_reg_b = "CLOCK0",
    altsyncram_component.indata_reg_b = "CLOCK0",
    altsyncram_component.wrcontrol_wraddress_reg_b = "CLOCK0",
    altsyncram_component.clock_enable_input_a = "BYPASS",
    altsyncram_component.clock_enable_output_a = "BYPASS",
    altsyncram_component.outdata_aclr_a = "NONE",
    altsyncram_component.outdata_reg_a = output_registered,
    altsyncram_component.numwords_a = numwords_a,
    altsyncram_component.widthad_a = widthad_a,
    altsyncram_component.width_a = width_a;

always @(*) begin
	clk_wire = clk;
end


endmodule
